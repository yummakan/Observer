LIBRARY ieee;
USE ieee.std_logic_1164.all;
use IEEE.NUMERIC_STD.ALL;

ENTITY TOP IS

PORT (

   clk 		:IN	std_logic;
	reset		:IN 	std_logic;
	
)

END TOP;
