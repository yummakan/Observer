LIBRARY ieee  ; 
LIBRARY std  ; 
USE ieee.NUMERIC_STD.all  ; 
USE ieee.std_logic_1164.all  ; 
USE ieee.std_logic_textio.all  ; 
USE ieee.std_logic_unsigned.all  ; 
USE std.textio.all  ; 
ENTITY \testbench_2.vhd\  IS 
END ; 
 
ARCHITECTURE \testbench_2.vhd_arch\   OF \testbench_2.vhd\   IS
  SIGNAL output   :  STD_LOGIC  ; 
  SIGNAL clk   :  STD_LOGIC  ; 
  SIGNAL reset   :  STD_LOGIC  ; 
  COMPONENT signalgenerator  
    PORT ( 
      output  : out STD_LOGIC ; 
      clk  : in STD_LOGIC ; 
      reset  : in STD_LOGIC ); 
  END COMPONENT ; 
BEGIN
  DUT  : signalgenerator 
    PORT MAP ( 
      output   => output  ,
      clk   => clk  ,
      reset   => reset   ) ; 



-- "Clock Pattern" : dutyCycle = 50
-- Start Time = 0 ns, End Time = 10 us, Period = 40 ns
  Process
	Begin
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
	 clk  <= '0'  ;
	wait for 20 ns ;
	 clk  <= '1'  ;
	wait for 20 ns ;
-- dumped values till 10 us
	wait;
 End Process;
 
 reset <= '1';
 
END;
